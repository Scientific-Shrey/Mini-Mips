`timescale 1ns/1ps

module register_file (
    input clk,
    input reg_write,
    input [4:0] read_reg1,
    input [4:0] read_reg2,
    input [4:0] write_reg,
    input [31:0] write_data,
    output [31:0] read_data1,
    output [31:0] read_data2
);
    reg [31:0] registers [0:31];//32 32 bit registers

    // Read operations
    assign read_data1 = registers[read_reg1];//read data
    assign read_data2 = registers[read_reg2];

    // Write operation
    always @(posedge clk) begin
        if (reg_write)//whenever reg_write, you write data
            registers[write_reg] <= write_data;
    end
endmodule
